library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PulseTimer is

	port(
		t_clear : in std_logic;
		sys_clk : in std_logic;
		dout	  : out std_logic_vector(9 downto 0)
	);

end entity;

architecture behaviour of PulseTimer is
	signal counter : integer;
begin

	process(sys_clk)
	begin
		if rising_edge(sys_clk) then
			if t_clear = '1' then
				counter <= 0 after 5 ns;
			else
				counter <= counter + 1 after 5 ns;
			end if;
		end if;
	end process;
	
	dout <= std_logic_vector(to_unsigned(counter,10));

end architecture;